module bft(
    input clk,
    input  [49-1:0]dout_leaf_0,
    input  [49-1:0]dout_leaf_1,
    input  [49-1:0]dout_leaf_2,
    input  [49-1:0]dout_leaf_3,
    input  [49-1:0]dout_leaf_4,
    input  [49-1:0]dout_leaf_5,
    input  [49-1:0]dout_leaf_6,
    input  [49-1:0]dout_leaf_7,
    input  [49-1:0]dout_leaf_8,
    input  [49-1:0]dout_leaf_9,
    input  [49-1:0]dout_leaf_10,
    input  [49-1:0]dout_leaf_11,
    input  [49-1:0]dout_leaf_12,
    input  [49-1:0]dout_leaf_13,
    input  [49-1:0]dout_leaf_14,
    input  [49-1:0]dout_leaf_15,
    output [49-1:0]din_leaf_0,
    output [49-1:0]din_leaf_1,
    output [49-1:0]din_leaf_2,
    output [49-1:0]din_leaf_3,
    output [49-1:0]din_leaf_4,
    output [49-1:0]din_leaf_5,
    output [49-1:0]din_leaf_6,
    output [49-1:0]din_leaf_7,
    output [49-1:0]din_leaf_8,
    output [49-1:0]din_leaf_9,
    output [49-1:0]din_leaf_10,
    output [49-1:0]din_leaf_11,
    output [49-1:0]din_leaf_12,
    output [49-1:0]din_leaf_13,
    output [49-1:0]din_leaf_14,
    output [49-1:0]din_leaf_15,
    output resend_0,
    output resend_1,
    output resend_2,
    output resend_3,
    output resend_4,
    output resend_5,
    output resend_6,
    output resend_7,
    output resend_8,
    output resend_9,
    output resend_10,
    output resend_11,
    output resend_12,
    output resend_13,
    output resend_14,
    output resend_15,
    input reset);
gen_nw16 # (        .num_leaves(16),
    .payload_sz(44),
    .p_sz(49),
    .addr(1'b0),
    .level(0)
    ) gen_nw16 (
    .clk(clk),
    .reset(reset),
    .pe_interface({
    dout_leaf_15,
    dout_leaf_14,
    dout_leaf_13,
    dout_leaf_12,
    dout_leaf_11,
    dout_leaf_10,
    dout_leaf_9,
    dout_leaf_8,
    dout_leaf_7,
    dout_leaf_6,
    dout_leaf_5,
    dout_leaf_4,
    dout_leaf_3,
    dout_leaf_2,
    dout_leaf_1,
    dout_leaf_0}),
    .interface_pe({
    din_leaf_15,
    din_leaf_14,
    din_leaf_13,
    din_leaf_12,
    din_leaf_11,
    din_leaf_10,
    din_leaf_9,
    din_leaf_8,
    din_leaf_7,
    din_leaf_6,
    din_leaf_5,
    din_leaf_4,
    din_leaf_3,
    din_leaf_2,
    din_leaf_1,
    din_leaf_0}),
    .resend({
    resend_15,
    resend_14,
    resend_13,
    resend_12,
    resend_11,
    resend_10,
    resend_9,
    resend_8,
    resend_7,
    resend_6,
    resend_5,
    resend_4,
    resend_3,
    resend_2,
    resend_1,
    resend_0}));
endmodule
